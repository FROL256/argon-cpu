 signal program  : PROGRAM_MEMORY  := 
 ( 
  0 => x"C1100000",
  1 => x"00000003",
  2 => x"C1200000",
  3 => x"00000002",
  4 => x"42012000",
  5 => x"12000000",
  6 => x"12000000",
  7 => x"12000000",
  others => x"00000000"
  );  
  
  
  
i, 1, a, mov, R1 
d, {3}
i, 1, a, mov, R2
d, {2}
r, 1, a, add, R0, R1, R2
r, 0, c, hlt, 0, 0, 0
r, 0, c, hlt, 0, 0, 0
r, 0, c, hlt, 0, 0, 0
